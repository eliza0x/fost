`include "../CPU.sv"
`include "../src/Parameter.sv"

module Add2();
    bit board_ck;
    bit CLK;
    bit rst;
    bit do_halt;
    logic [7:0] SEG_A,SEG_B,SEG_C,SEG_D,SEG_E,SEG_F,SEG_G,SEG_H;
    logic [8:0] SEG_SEL_IK;
    logic [7:0] SEG;
    logic [3:0] SEG_SEL;

    CPU cpu(.*);

    always #(one_clock*2) board_ck = ~board_ck;

    always @(negedge do_halt) begin
        $display("=================================");
        for (byte i=0; i<10; i++) begin
            $display("memory[%2d]: %d", i, cpu.memory_module.memory[i]);
        end
        $display("--------------------------------");
        for (byte i=0; i<16; i++) begin
            $display("regs[%2d]: %d", i, cpu.decode_module.regs[i]);
        end
        $display("=================================");

        $display("regs[1]: %d", cpu.decode_module.regs[1]);
        $display("regs[2]: %d", cpu.decode_module.regs[2]);
        assert(cpu.decode_module.regs[1] == 12);
        assert(cpu.decode_module.regs[2] == 5);

        $finish(1);
    end

    initial begin
        $display("do_halt: %d", do_halt);
        board_ck = 1'b0;
        rst = 1;

        cpu.fetch_module.memory[ 0] <= 16'h0000;
        cpu.fetch_module.memory[ 1] <= 16'b1000_0001_00000111 ; // ldi
        cpu.fetch_module.memory[ 2] <= 16'b1000_0010_00000101 ; // ldi
        cpu.fetch_module.memory[ 3] <= 16'b0001_0001_0010_0000; // add 
        cpu.fetch_module.memory[ 4] <= 16'b1111111111111111   ; // halt

        #100000 $finish(1);
    end
endmodule
