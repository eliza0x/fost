// 動作周波数
parameter one_clock = 50;

parameter op_begin = 15;
parameter op_end   = 12;

parameter rd_begin = 11;
parameter rd_end   = 8;

parameter rs_begin = 7;
parameter rs_end   = 4;

parameter rt_begin = 3;
parameter rt_end   = 0;

parameter i9_begin = 8;
parameter i9_end   = 0;

